module my_module(input r1, input r2, output c, output d);
add r1, r2, r3
if (r1 == r2) r3 = r1 + r2;
for (i = 0; i < 10; i = i + 1) begin
endmodule